library IEEE;
use ieee.std_logic_1164.all;

entity morse_code_encoder is
	port ();
end morse_code_encoder;
